* Super simple RC test circuit
V1 VIN 0 0 AC 1 0
R1 VOUT VIN 1k
C1 VOUT 0 159n
.ac dec 10 1 1Meg
.plot ac VOUT
.end