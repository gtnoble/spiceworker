* MOSFET RF Amplifier objective function

.SUBCKT irf510 1 2 3
* Model generated on Apr 24, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=3.82703 LAMBDA=0 KP=2.48457
+CGSO=1.72132e-06 CGDO=5.99235e-11
RS 8 3 0.276929
D1 3 1 MD
.MODEL MD D IS=6.52734e-11 RS=0.0458243 N=1.2565 BV=100
+IBV=0.00025 EG=1.2 XTI=1 TT=0
+CJO=2.98645e-10 VJ=0.774158 M=0.422859 FC=0.5
RDS 3 1 4e+06
RD 9 1 0.0673242
RG 2 7 13.1694
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.85121e-10 VJ=0.500044 M=0.651006 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.40332e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS

XMOS1 N010 N011 N012 IRF510
L§INPUT_CHOKE N008 N015 1m
L§OUTPUT_CHOKE V+ N001 1m
V1 V+ 0 12
V2 VIN 0 0 AC 10m
R§INPUT_IMPEDANCE N013 VIN 50
R§SOURCE_RESISTOR N017 0 0.219561254573105
C§OUTPUT_DC_BLOCK N002 N001 8.16120626212353e-05
R§OUTPUT_IMPEDANCE VOUT 0 50
L§GATE_PARASITIC_L N016 N015 5n
R§GATE_PARASITIC_R N011 N016 30m
L§SOURCE_PARASITIC_L N012 N017 5n
L§DRAIN_PARASITIC_L N009 N010 1.88n
L§INPUT_SECONDARY N014 0 4.9988835944874e-05
L§INPUT_PRIMARY N013 0 0.000223162548486584
L§OUTPUT_PRIMARY N002 0 3.71525795216264e-05
L§OUTPUT_SECONDARY VOUT 0 9.45258187936205e-05
XMOS2 N005 N006 N007 IRF510
R§GATE_PARASITIC_R1 N006 N004 30m
L§SOURCE_PARASITIC_L1 N007 N009 5n
L§DRAIN_PARASITIC_L1 N001 N005 1.88n
C§SECONDARY_DC_BLOCK N015 N014 1.27723941412898e-05
V§COMMON_GATE_BIAS N003 0 9.08849117036013
V§EMITTER_FOLLOWER_BIAS N008 0 4.26815040170132
L§GATE_PARASITIC_L1 N004 N003 5n

KOUTPUT L§OUTPUT_PRIMARY L§OUTPUT_SECONDARY 1
KINPUT L§INPUT_PRIMARY L§INPUT_SECONDARY 1

.probe p(XMOS1)
.probe p(XMOS2)

.op
.control
  run

  let objective = (vecmin(mag(VOUT)))

  wrdata $tempFile objective
  quit
.endc

.end


